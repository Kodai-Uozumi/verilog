library verilog;
use verilog.vl_types.all;
entity adder2_test is
    generic(
        STEP            : integer := 1000
    );
end adder2_test;
