library verilog;
use verilog.vl_types.all;
entity prienc_test is
    generic(
        STEP            : integer := 1000
    );
end prienc_test;
