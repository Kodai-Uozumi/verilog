library verilog;
use verilog.vl_types.all;
entity up256_test is
    generic(
        STEP            : integer := 1000
    );
end up256_test;
