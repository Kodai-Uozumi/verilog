library verilog;
use verilog.vl_types.all;
entity down3_test is
    generic(
        STEP            : integer := 1000
    );
end down3_test;
