library verilog;
use verilog.vl_types.all;
entity comp2_test is
    generic(
        STEP            : integer := 1000
    );
end comp2_test;
