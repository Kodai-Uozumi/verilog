library verilog;
use verilog.vl_types.all;
entity up4_test is
    generic(
        STEP            : integer := 1000
    );
end up4_test;
